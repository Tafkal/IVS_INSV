-- system.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk       : in    std_logic                     := '0';             --       clk.clk
		reset_reset_n : in    std_logic                     := '0';             --     reset.reset_n
		sdram_addr    : out   std_logic_vector(11 downto 0);                    --     sdram.addr
		sdram_ba      : out   std_logic_vector(1 downto 0);                     --          .ba
		sdram_cas_n   : out   std_logic;                                        --          .cas_n
		sdram_cke     : out   std_logic;                                        --          .cke
		sdram_cs_n    : out   std_logic;                                        --          .cs_n
		sdram_dq      : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		sdram_dqm     : out   std_logic_vector(1 downto 0);                     --          .dqm
		sdram_ras_n   : out   std_logic;                                        --          .ras_n
		sdram_we_n    : out   std_logic;                                        --          .we_n
		sdram_clk_clk : out   std_logic                                         -- sdram_clk.clk
	);
end entity system;

architecture rtl of system is
	component system_ack_fifo is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			wrreset_n                        : in  std_logic                     := 'X';             -- reset_n
			rdclock                          : in  std_logic                     := 'X';             -- clk
			rdreset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			rdclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			rdclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			rdclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rdclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			rdclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component system_ack_fifo;

	component system_manager is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_manager;

	component system_manager_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_manager_jtag_uart;

	component system_mutex is
		port (
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk           : in  std_logic                     := 'X';             -- clk
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			address       : in  std_logic                     := 'X'              -- address
		);
	end component system_mutex;

	component system_pcu is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component system_pcu;

	component system_pll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component system_pll_0;

	component system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_sdram;

	component system_shared_ocm is
		port (
			address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component system_shared_ocm;

	component system_workers is
		port (
			clk_clk            : in  std_logic                     := 'X';             -- clk
			reset_reset_n      : in  std_logic                     := 'X';             -- reset_n
			wout_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			wout_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			wout_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			wout_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			wout_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			wout_address       : out std_logic_vector(27 downto 0);                    -- address
			wout_write         : out std_logic;                                        -- write
			wout_read          : out std_logic;                                        -- read
			wout_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			wout_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component system_workers;

	component system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			pll_0_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			manager_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			pll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			workers_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			manager_data_master_address                             : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			manager_data_master_waitrequest                         : out std_logic;                                        -- waitrequest
			manager_data_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			manager_data_master_read                                : in  std_logic                     := 'X';             -- read
			manager_data_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			manager_data_master_readdatavalid                       : out std_logic;                                        -- readdatavalid
			manager_data_master_write                               : in  std_logic                     := 'X';             -- write
			manager_data_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			manager_data_master_debugaccess                         : in  std_logic                     := 'X';             -- debugaccess
			manager_instruction_master_address                      : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			manager_instruction_master_waitrequest                  : out std_logic;                                        -- waitrequest
			manager_instruction_master_read                         : in  std_logic                     := 'X';             -- read
			manager_instruction_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			manager_instruction_master_readdatavalid                : out std_logic;                                        -- readdatavalid
			workers_wout_address                                    : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			workers_wout_waitrequest                                : out std_logic;                                        -- waitrequest
			workers_wout_burstcount                                 : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			workers_wout_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			workers_wout_read                                       : in  std_logic                     := 'X';             -- read
			workers_wout_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			workers_wout_readdatavalid                              : out std_logic;                                        -- readdatavalid
			workers_wout_write                                      : in  std_logic                     := 'X';             -- write
			workers_wout_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			workers_wout_debugaccess                                : in  std_logic                     := 'X';             -- debugaccess
			ack_fifo_in_write                                       : out std_logic;                                        -- write
			ack_fifo_in_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			ack_fifo_in_waitrequest                                 : in  std_logic                     := 'X';             -- waitrequest
			ack_fifo_in_csr_address                                 : out std_logic_vector(2 downto 0);                     -- address
			ack_fifo_in_csr_write                                   : out std_logic;                                        -- write
			ack_fifo_in_csr_read                                    : out std_logic;                                        -- read
			ack_fifo_in_csr_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ack_fifo_in_csr_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			ack_fifo_out_read                                       : out std_logic;                                        -- read
			ack_fifo_out_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ack_fifo_out_waitrequest                                : in  std_logic                     := 'X';             -- waitrequest
			ack_fifo_out_csr_address                                : out std_logic_vector(2 downto 0);                     -- address
			ack_fifo_out_csr_write                                  : out std_logic;                                        -- write
			ack_fifo_out_csr_read                                   : out std_logic;                                        -- read
			ack_fifo_out_csr_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ack_fifo_out_csr_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			manager_debug_mem_slave_address                         : out std_logic_vector(8 downto 0);                     -- address
			manager_debug_mem_slave_write                           : out std_logic;                                        -- write
			manager_debug_mem_slave_read                            : out std_logic;                                        -- read
			manager_debug_mem_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			manager_debug_mem_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			manager_debug_mem_slave_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			manager_debug_mem_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			manager_debug_mem_slave_debugaccess                     : out std_logic;                                        -- debugaccess
			manager_jtag_uart_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			manager_jtag_uart_avalon_jtag_slave_write               : out std_logic;                                        -- write
			manager_jtag_uart_avalon_jtag_slave_read                : out std_logic;                                        -- read
			manager_jtag_uart_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			manager_jtag_uart_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			manager_jtag_uart_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			manager_jtag_uart_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			mutex_s1_address                                        : out std_logic_vector(0 downto 0);                     -- address
			mutex_s1_write                                          : out std_logic;                                        -- write
			mutex_s1_read                                           : out std_logic;                                        -- read
			mutex_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mutex_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			mutex_s1_chipselect                                     : out std_logic;                                        -- chipselect
			pcu_control_slave_address                               : out std_logic_vector(2 downto 0);                     -- address
			pcu_control_slave_write                                 : out std_logic;                                        -- write
			pcu_control_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pcu_control_slave_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pcu_control_slave_begintransfer                         : out std_logic;                                        -- begintransfer
			pll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_0_pll_slave_write                                   : out std_logic;                                        -- write
			pll_0_pll_slave_read                                    : out std_logic;                                        -- read
			pll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_s1_address                                        : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                                          : out std_logic;                                        -- write
			sdram_s1_read                                           : out std_logic;                                        -- read
			sdram_s1_readdata                                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                      : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                     : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                     : out std_logic;                                        -- chipselect
			shared_ocm_s1_address                                   : out std_logic_vector(7 downto 0);                     -- address
			shared_ocm_s1_write                                     : out std_logic;                                        -- write
			shared_ocm_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			shared_ocm_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			shared_ocm_s1_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			shared_ocm_s1_chipselect                                : out std_logic;                                        -- chipselect
			shared_ocm_s1_clken                                     : out std_logic;                                        -- clken
			shared_ocm_s2_address                                   : out std_logic_vector(7 downto 0);                     -- address
			shared_ocm_s2_write                                     : out std_logic;                                        -- write
			shared_ocm_s2_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			shared_ocm_s2_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			shared_ocm_s2_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			shared_ocm_s2_chipselect                                : out std_logic;                                        -- chipselect
			shared_ocm_s2_clken                                     : out std_logic                                         -- clken
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	signal pll_0_c0_clk                                                          : std_logic;                     -- pll_0:c0 -> [ack_fifo:rdclock, ack_fifo:wrclock, irq_mapper:clk, manager:clk, manager_jtag_uart:clk, mm_interconnect_0:pll_0_c0_clk, mutex:clk, pcu:clk, rst_controller:clk, sdram:clk, shared_ocm:clk, workers:clk_clk]
	signal manager_data_master_readdata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_data_master_readdata -> manager:d_readdata
	signal manager_data_master_waitrequest                                       : std_logic;                     -- mm_interconnect_0:manager_data_master_waitrequest -> manager:d_waitrequest
	signal manager_data_master_debugaccess                                       : std_logic;                     -- manager:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:manager_data_master_debugaccess
	signal manager_data_master_address                                           : std_logic_vector(26 downto 0); -- manager:d_address -> mm_interconnect_0:manager_data_master_address
	signal manager_data_master_byteenable                                        : std_logic_vector(3 downto 0);  -- manager:d_byteenable -> mm_interconnect_0:manager_data_master_byteenable
	signal manager_data_master_read                                              : std_logic;                     -- manager:d_read -> mm_interconnect_0:manager_data_master_read
	signal manager_data_master_readdatavalid                                     : std_logic;                     -- mm_interconnect_0:manager_data_master_readdatavalid -> manager:d_readdatavalid
	signal manager_data_master_write                                             : std_logic;                     -- manager:d_write -> mm_interconnect_0:manager_data_master_write
	signal manager_data_master_writedata                                         : std_logic_vector(31 downto 0); -- manager:d_writedata -> mm_interconnect_0:manager_data_master_writedata
	signal manager_instruction_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_instruction_master_readdata -> manager:i_readdata
	signal manager_instruction_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:manager_instruction_master_waitrequest -> manager:i_waitrequest
	signal manager_instruction_master_address                                    : std_logic_vector(26 downto 0); -- manager:i_address -> mm_interconnect_0:manager_instruction_master_address
	signal manager_instruction_master_read                                       : std_logic;                     -- manager:i_read -> mm_interconnect_0:manager_instruction_master_read
	signal manager_instruction_master_readdatavalid                              : std_logic;                     -- mm_interconnect_0:manager_instruction_master_readdatavalid -> manager:i_readdatavalid
	signal workers_wout_waitrequest                                              : std_logic;                     -- mm_interconnect_0:workers_wout_waitrequest -> workers:wout_waitrequest
	signal workers_wout_readdata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:workers_wout_readdata -> workers:wout_readdata
	signal workers_wout_debugaccess                                              : std_logic;                     -- workers:wout_debugaccess -> mm_interconnect_0:workers_wout_debugaccess
	signal workers_wout_address                                                  : std_logic_vector(27 downto 0); -- workers:wout_address -> mm_interconnect_0:workers_wout_address
	signal workers_wout_read                                                     : std_logic;                     -- workers:wout_read -> mm_interconnect_0:workers_wout_read
	signal workers_wout_byteenable                                               : std_logic_vector(3 downto 0);  -- workers:wout_byteenable -> mm_interconnect_0:workers_wout_byteenable
	signal workers_wout_readdatavalid                                            : std_logic;                     -- mm_interconnect_0:workers_wout_readdatavalid -> workers:wout_readdatavalid
	signal workers_wout_writedata                                                : std_logic_vector(31 downto 0); -- workers:wout_writedata -> mm_interconnect_0:workers_wout_writedata
	signal workers_wout_write                                                    : std_logic;                     -- workers:wout_write -> mm_interconnect_0:workers_wout_write
	signal workers_wout_burstcount                                               : std_logic_vector(0 downto 0);  -- workers:wout_burstcount -> mm_interconnect_0:workers_wout_burstcount
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_chipselect -> manager_jtag_uart:av_chipselect
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- manager_jtag_uart:av_readdata -> mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- manager_jtag_uart:av_waitrequest -> mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_address -> manager_jtag_uart:av_address
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_writedata -> manager_jtag_uart:av_writedata
	signal mm_interconnect_0_pcu_control_slave_readdata                          : std_logic_vector(31 downto 0); -- pcu:readdata -> mm_interconnect_0:pcu_control_slave_readdata
	signal mm_interconnect_0_pcu_control_slave_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pcu_control_slave_address -> pcu:address
	signal mm_interconnect_0_pcu_control_slave_begintransfer                     : std_logic;                     -- mm_interconnect_0:pcu_control_slave_begintransfer -> pcu:begintransfer
	signal mm_interconnect_0_pcu_control_slave_write                             : std_logic;                     -- mm_interconnect_0:pcu_control_slave_write -> pcu:write
	signal mm_interconnect_0_pcu_control_slave_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:pcu_control_slave_writedata -> pcu:writedata
	signal mm_interconnect_0_manager_debug_mem_slave_readdata                    : std_logic_vector(31 downto 0); -- manager:debug_mem_slave_readdata -> mm_interconnect_0:manager_debug_mem_slave_readdata
	signal mm_interconnect_0_manager_debug_mem_slave_waitrequest                 : std_logic;                     -- manager:debug_mem_slave_waitrequest -> mm_interconnect_0:manager_debug_mem_slave_waitrequest
	signal mm_interconnect_0_manager_debug_mem_slave_debugaccess                 : std_logic;                     -- mm_interconnect_0:manager_debug_mem_slave_debugaccess -> manager:debug_mem_slave_debugaccess
	signal mm_interconnect_0_manager_debug_mem_slave_address                     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:manager_debug_mem_slave_address -> manager:debug_mem_slave_address
	signal mm_interconnect_0_manager_debug_mem_slave_read                        : std_logic;                     -- mm_interconnect_0:manager_debug_mem_slave_read -> manager:debug_mem_slave_read
	signal mm_interconnect_0_manager_debug_mem_slave_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:manager_debug_mem_slave_byteenable -> manager:debug_mem_slave_byteenable
	signal mm_interconnect_0_manager_debug_mem_slave_write                       : std_logic;                     -- mm_interconnect_0:manager_debug_mem_slave_write -> manager:debug_mem_slave_write
	signal mm_interconnect_0_manager_debug_mem_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_debug_mem_slave_writedata -> manager:debug_mem_slave_writedata
	signal mm_interconnect_0_ack_fifo_out_readdata                               : std_logic_vector(31 downto 0); -- ack_fifo:avalonmm_read_slave_readdata -> mm_interconnect_0:ack_fifo_out_readdata
	signal mm_interconnect_0_ack_fifo_out_waitrequest                            : std_logic;                     -- ack_fifo:avalonmm_read_slave_waitrequest -> mm_interconnect_0:ack_fifo_out_waitrequest
	signal mm_interconnect_0_ack_fifo_out_read                                   : std_logic;                     -- mm_interconnect_0:ack_fifo_out_read -> ack_fifo:avalonmm_read_slave_read
	signal mm_interconnect_0_ack_fifo_out_csr_readdata                           : std_logic_vector(31 downto 0); -- ack_fifo:rdclk_control_slave_readdata -> mm_interconnect_0:ack_fifo_out_csr_readdata
	signal mm_interconnect_0_ack_fifo_out_csr_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ack_fifo_out_csr_address -> ack_fifo:rdclk_control_slave_address
	signal mm_interconnect_0_ack_fifo_out_csr_read                               : std_logic;                     -- mm_interconnect_0:ack_fifo_out_csr_read -> ack_fifo:rdclk_control_slave_read
	signal mm_interconnect_0_ack_fifo_out_csr_write                              : std_logic;                     -- mm_interconnect_0:ack_fifo_out_csr_write -> ack_fifo:rdclk_control_slave_write
	signal mm_interconnect_0_ack_fifo_out_csr_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:ack_fifo_out_csr_writedata -> ack_fifo:rdclk_control_slave_writedata
	signal mm_interconnect_0_pll_0_pll_slave_readdata                            : std_logic_vector(31 downto 0); -- pll_0:readdata -> mm_interconnect_0:pll_0_pll_slave_readdata
	signal mm_interconnect_0_pll_0_pll_slave_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_0_pll_slave_address -> pll_0:address
	signal mm_interconnect_0_pll_0_pll_slave_read                                : std_logic;                     -- mm_interconnect_0:pll_0_pll_slave_read -> pll_0:read
	signal mm_interconnect_0_pll_0_pll_slave_write                               : std_logic;                     -- mm_interconnect_0:pll_0_pll_slave_write -> pll_0:write
	signal mm_interconnect_0_pll_0_pll_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_0_pll_slave_writedata -> pll_0:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                   : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                    : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                       : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                              : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                      : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_shared_ocm_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:shared_ocm_s1_chipselect -> shared_ocm:chipselect
	signal mm_interconnect_0_shared_ocm_s1_readdata                              : std_logic_vector(31 downto 0); -- shared_ocm:readdata -> mm_interconnect_0:shared_ocm_s1_readdata
	signal mm_interconnect_0_shared_ocm_s1_address                               : std_logic_vector(7 downto 0);  -- mm_interconnect_0:shared_ocm_s1_address -> shared_ocm:address
	signal mm_interconnect_0_shared_ocm_s1_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:shared_ocm_s1_byteenable -> shared_ocm:byteenable
	signal mm_interconnect_0_shared_ocm_s1_write                                 : std_logic;                     -- mm_interconnect_0:shared_ocm_s1_write -> shared_ocm:write
	signal mm_interconnect_0_shared_ocm_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:shared_ocm_s1_writedata -> shared_ocm:writedata
	signal mm_interconnect_0_shared_ocm_s1_clken                                 : std_logic;                     -- mm_interconnect_0:shared_ocm_s1_clken -> shared_ocm:clken
	signal mm_interconnect_0_mutex_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:mutex_s1_chipselect -> mutex:chipselect
	signal mm_interconnect_0_mutex_s1_readdata                                   : std_logic_vector(31 downto 0); -- mutex:data_to_cpu -> mm_interconnect_0:mutex_s1_readdata
	signal mm_interconnect_0_mutex_s1_address                                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mutex_s1_address -> mutex:address
	signal mm_interconnect_0_mutex_s1_read                                       : std_logic;                     -- mm_interconnect_0:mutex_s1_read -> mutex:read
	signal mm_interconnect_0_mutex_s1_write                                      : std_logic;                     -- mm_interconnect_0:mutex_s1_write -> mutex:write
	signal mm_interconnect_0_mutex_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:mutex_s1_writedata -> mutex:data_from_cpu
	signal mm_interconnect_0_ack_fifo_in_waitrequest                             : std_logic;                     -- ack_fifo:avalonmm_write_slave_waitrequest -> mm_interconnect_0:ack_fifo_in_waitrequest
	signal mm_interconnect_0_ack_fifo_in_write                                   : std_logic;                     -- mm_interconnect_0:ack_fifo_in_write -> ack_fifo:avalonmm_write_slave_write
	signal mm_interconnect_0_ack_fifo_in_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:ack_fifo_in_writedata -> ack_fifo:avalonmm_write_slave_writedata
	signal mm_interconnect_0_ack_fifo_in_csr_readdata                            : std_logic_vector(31 downto 0); -- ack_fifo:wrclk_control_slave_readdata -> mm_interconnect_0:ack_fifo_in_csr_readdata
	signal mm_interconnect_0_ack_fifo_in_csr_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ack_fifo_in_csr_address -> ack_fifo:wrclk_control_slave_address
	signal mm_interconnect_0_ack_fifo_in_csr_read                                : std_logic;                     -- mm_interconnect_0:ack_fifo_in_csr_read -> ack_fifo:wrclk_control_slave_read
	signal mm_interconnect_0_ack_fifo_in_csr_write                               : std_logic;                     -- mm_interconnect_0:ack_fifo_in_csr_write -> ack_fifo:wrclk_control_slave_write
	signal mm_interconnect_0_ack_fifo_in_csr_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:ack_fifo_in_csr_writedata -> ack_fifo:wrclk_control_slave_writedata
	signal mm_interconnect_0_shared_ocm_s2_chipselect                            : std_logic;                     -- mm_interconnect_0:shared_ocm_s2_chipselect -> shared_ocm:chipselect2
	signal mm_interconnect_0_shared_ocm_s2_readdata                              : std_logic_vector(31 downto 0); -- shared_ocm:readdata2 -> mm_interconnect_0:shared_ocm_s2_readdata
	signal mm_interconnect_0_shared_ocm_s2_address                               : std_logic_vector(7 downto 0);  -- mm_interconnect_0:shared_ocm_s2_address -> shared_ocm:address2
	signal mm_interconnect_0_shared_ocm_s2_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:shared_ocm_s2_byteenable -> shared_ocm:byteenable2
	signal mm_interconnect_0_shared_ocm_s2_write                                 : std_logic;                     -- mm_interconnect_0:shared_ocm_s2_write -> shared_ocm:write2
	signal mm_interconnect_0_shared_ocm_s2_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:shared_ocm_s2_writedata -> shared_ocm:writedata2
	signal mm_interconnect_0_shared_ocm_s2_clken                                 : std_logic;                     -- mm_interconnect_0:shared_ocm_s2_clken -> shared_ocm:clken2
	signal irq_mapper_receiver0_irq                                              : std_logic;                     -- manager_jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal manager_irq_irq                                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> manager:irq
	signal rst_controller_reset_out_reset                                        : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:manager_reset_reset_bridge_in_reset_reset, mm_interconnect_0:workers_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, shared_ocm:reset]
	signal rst_controller_reset_out_reset_req                                    : std_logic;                     -- rst_controller:reset_req -> [manager:reset_req, rst_translator:reset_req_in, shared_ocm:reset_req]
	signal manager_debug_reset_request_reset                                     : std_logic;                     -- manager:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                                    : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pll_0_inclk_interface_reset_reset_bridge_in_reset_reset, pll_0:reset]
	signal rst_controller_002_reset_out_reset                                    : std_logic;                     -- rst_controller_002:reset_out -> rst_controller_002_reset_out_reset:in
	signal reset_reset_n_ports_inv                                               : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read:inv -> manager_jtag_uart:av_read_n
	signal mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write:inv -> manager_jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                             : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_reset_out_reset:inv -> [ack_fifo:rdreset_n, ack_fifo:wrreset_n, manager:reset_n, manager_jtag_uart:rst_n, mutex:reset_n, pcu:reset_n, sdram:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> workers:reset_reset_n

begin

	ack_fifo : component system_ack_fifo
		port map (
			wrclock                          => pll_0_c0_clk,                                 --    clk_in.clk
			wrreset_n                        => rst_controller_reset_out_reset_ports_inv,     --  reset_in.reset_n
			rdclock                          => pll_0_c0_clk,                                 --   clk_out.clk
			rdreset_n                        => rst_controller_reset_out_reset_ports_inv,     -- reset_out.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_0_ack_fifo_in_writedata,      --        in.writedata
			avalonmm_write_slave_write       => mm_interconnect_0_ack_fifo_in_write,          --          .write
			avalonmm_write_slave_waitrequest => mm_interconnect_0_ack_fifo_in_waitrequest,    --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_0_ack_fifo_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_0_ack_fifo_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_0_ack_fifo_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_0_ack_fifo_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_0_ack_fifo_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_0_ack_fifo_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_0_ack_fifo_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_0_ack_fifo_out_csr_readdata,  --          .readdata
			wrclk_control_slave_address      => mm_interconnect_0_ack_fifo_in_csr_address,    --    in_csr.address
			wrclk_control_slave_read         => mm_interconnect_0_ack_fifo_in_csr_read,       --          .read
			wrclk_control_slave_writedata    => mm_interconnect_0_ack_fifo_in_csr_writedata,  --          .writedata
			wrclk_control_slave_write        => mm_interconnect_0_ack_fifo_in_csr_write,      --          .write
			wrclk_control_slave_readdata     => mm_interconnect_0_ack_fifo_in_csr_readdata    --          .readdata
		);

	manager : component system_manager
		port map (
			clk                                 => pll_0_c0_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,              --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                           => manager_data_master_address,                           --               data_master.address
			d_byteenable                        => manager_data_master_byteenable,                        --                          .byteenable
			d_read                              => manager_data_master_read,                              --                          .read
			d_readdata                          => manager_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => manager_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => manager_data_master_write,                             --                          .write
			d_writedata                         => manager_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => manager_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => manager_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => manager_instruction_master_address,                    --        instruction_master.address
			i_read                              => manager_instruction_master_read,                       --                          .read
			i_readdata                          => manager_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => manager_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => manager_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => manager_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => manager_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_manager_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_manager_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_manager_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_manager_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_manager_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_manager_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_manager_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_manager_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	manager_jtag_uart : component system_manager_jtag_uart
		port map (
			clk            => pll_0_c0_clk,                                                          --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                              --             reset.reset_n
			av_chipselect  => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                               --               irq.irq
		);

	mutex : component system_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv, -- reset.reset_n
			clk           => pll_0_c0_clk,                             --   clk.clk
			chipselect    => mm_interconnect_0_mutex_s1_chipselect,    --    s1.chipselect
			data_from_cpu => mm_interconnect_0_mutex_s1_writedata,     --      .writedata
			read          => mm_interconnect_0_mutex_s1_read,          --      .read
			write         => mm_interconnect_0_mutex_s1_write,         --      .write
			data_to_cpu   => mm_interconnect_0_mutex_s1_readdata,      --      .readdata
			address       => mm_interconnect_0_mutex_s1_address(0)     --      .address
		);

	pcu : component system_pcu
		port map (
			clk           => pll_0_c0_clk,                                      --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			address       => mm_interconnect_0_pcu_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_pcu_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_pcu_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_pcu_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_pcu_control_slave_writedata      --              .writedata
		);

	pll_0 : component system_pll_0
		port map (
			clk                => clk_clk,                                     --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,          -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_0_pll_slave_writedata, --                      .writedata
			c0                 => pll_0_c0_clk,                                --                    c0.clk
			c1                 => sdram_clk_clk,                               --                    c1.clk
			scandone           => open,                                        --           (terminated)
			scandataout        => open,                                        --           (terminated)
			areset             => '0',                                         --           (terminated)
			locked             => open,                                        --           (terminated)
			phasedone          => open,                                        --           (terminated)
			phasecounterselect => "0000",                                      --           (terminated)
			phaseupdown        => '0',                                         --           (terminated)
			phasestep          => '0',                                         --           (terminated)
			scanclk            => '0',                                         --           (terminated)
			scanclkena         => '0',                                         --           (terminated)
			scandata           => '0',                                         --           (terminated)
			configupdate       => '0'                                          --           (terminated)
		);

	sdram : component system_sdram
		port map (
			clk            => pll_0_c0_clk,                                    --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	shared_ocm : component system_shared_ocm
		port map (
			address     => mm_interconnect_0_shared_ocm_s1_address,    --     s1.address
			clken       => mm_interconnect_0_shared_ocm_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_shared_ocm_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_shared_ocm_s1_write,      --       .write
			readdata    => mm_interconnect_0_shared_ocm_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_shared_ocm_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_shared_ocm_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_0_shared_ocm_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_shared_ocm_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_shared_ocm_s2_clken,      --       .clken
			write2      => mm_interconnect_0_shared_ocm_s2_write,      --       .write
			readdata2   => mm_interconnect_0_shared_ocm_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_shared_ocm_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_shared_ocm_s2_byteenable, --       .byteenable
			clk         => pll_0_c0_clk,                               --   clk1.clk
			reset       => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze      => '0'                                         -- (terminated)
		);

	workers : component system_workers
		port map (
			clk_clk            => pll_0_c0_clk,                                 --   clk.clk
			reset_reset_n      => rst_controller_002_reset_out_reset_ports_inv, -- reset.reset_n
			wout_waitrequest   => workers_wout_waitrequest,                     --  wout.waitrequest
			wout_readdata      => workers_wout_readdata,                        --      .readdata
			wout_readdatavalid => workers_wout_readdatavalid,                   --      .readdatavalid
			wout_burstcount    => workers_wout_burstcount,                      --      .burstcount
			wout_writedata     => workers_wout_writedata,                       --      .writedata
			wout_address       => workers_wout_address,                         --      .address
			wout_write         => workers_wout_write,                           --      .write
			wout_read          => workers_wout_read,                            --      .read
			wout_byteenable    => workers_wout_byteenable,                      --      .byteenable
			wout_debugaccess   => workers_wout_debugaccess                      --      .debugaccess
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                           => clk_clk,                                                           --                                         clk_0_clk.clk
			pll_0_c0_clk                                            => pll_0_c0_clk,                                                      --                                          pll_0_c0.clk
			manager_reset_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,                                    --               manager_reset_reset_bridge_in_reset.reset
			pll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                -- pll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			workers_reset_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,                                    --               workers_reset_reset_bridge_in_reset.reset
			manager_data_master_address                             => manager_data_master_address,                                       --                               manager_data_master.address
			manager_data_master_waitrequest                         => manager_data_master_waitrequest,                                   --                                                  .waitrequest
			manager_data_master_byteenable                          => manager_data_master_byteenable,                                    --                                                  .byteenable
			manager_data_master_read                                => manager_data_master_read,                                          --                                                  .read
			manager_data_master_readdata                            => manager_data_master_readdata,                                      --                                                  .readdata
			manager_data_master_readdatavalid                       => manager_data_master_readdatavalid,                                 --                                                  .readdatavalid
			manager_data_master_write                               => manager_data_master_write,                                         --                                                  .write
			manager_data_master_writedata                           => manager_data_master_writedata,                                     --                                                  .writedata
			manager_data_master_debugaccess                         => manager_data_master_debugaccess,                                   --                                                  .debugaccess
			manager_instruction_master_address                      => manager_instruction_master_address,                                --                        manager_instruction_master.address
			manager_instruction_master_waitrequest                  => manager_instruction_master_waitrequest,                            --                                                  .waitrequest
			manager_instruction_master_read                         => manager_instruction_master_read,                                   --                                                  .read
			manager_instruction_master_readdata                     => manager_instruction_master_readdata,                               --                                                  .readdata
			manager_instruction_master_readdatavalid                => manager_instruction_master_readdatavalid,                          --                                                  .readdatavalid
			workers_wout_address                                    => workers_wout_address,                                              --                                      workers_wout.address
			workers_wout_waitrequest                                => workers_wout_waitrequest,                                          --                                                  .waitrequest
			workers_wout_burstcount                                 => workers_wout_burstcount,                                           --                                                  .burstcount
			workers_wout_byteenable                                 => workers_wout_byteenable,                                           --                                                  .byteenable
			workers_wout_read                                       => workers_wout_read,                                                 --                                                  .read
			workers_wout_readdata                                   => workers_wout_readdata,                                             --                                                  .readdata
			workers_wout_readdatavalid                              => workers_wout_readdatavalid,                                        --                                                  .readdatavalid
			workers_wout_write                                      => workers_wout_write,                                                --                                                  .write
			workers_wout_writedata                                  => workers_wout_writedata,                                            --                                                  .writedata
			workers_wout_debugaccess                                => workers_wout_debugaccess,                                          --                                                  .debugaccess
			ack_fifo_in_write                                       => mm_interconnect_0_ack_fifo_in_write,                               --                                       ack_fifo_in.write
			ack_fifo_in_writedata                                   => mm_interconnect_0_ack_fifo_in_writedata,                           --                                                  .writedata
			ack_fifo_in_waitrequest                                 => mm_interconnect_0_ack_fifo_in_waitrequest,                         --                                                  .waitrequest
			ack_fifo_in_csr_address                                 => mm_interconnect_0_ack_fifo_in_csr_address,                         --                                   ack_fifo_in_csr.address
			ack_fifo_in_csr_write                                   => mm_interconnect_0_ack_fifo_in_csr_write,                           --                                                  .write
			ack_fifo_in_csr_read                                    => mm_interconnect_0_ack_fifo_in_csr_read,                            --                                                  .read
			ack_fifo_in_csr_readdata                                => mm_interconnect_0_ack_fifo_in_csr_readdata,                        --                                                  .readdata
			ack_fifo_in_csr_writedata                               => mm_interconnect_0_ack_fifo_in_csr_writedata,                       --                                                  .writedata
			ack_fifo_out_read                                       => mm_interconnect_0_ack_fifo_out_read,                               --                                      ack_fifo_out.read
			ack_fifo_out_readdata                                   => mm_interconnect_0_ack_fifo_out_readdata,                           --                                                  .readdata
			ack_fifo_out_waitrequest                                => mm_interconnect_0_ack_fifo_out_waitrequest,                        --                                                  .waitrequest
			ack_fifo_out_csr_address                                => mm_interconnect_0_ack_fifo_out_csr_address,                        --                                  ack_fifo_out_csr.address
			ack_fifo_out_csr_write                                  => mm_interconnect_0_ack_fifo_out_csr_write,                          --                                                  .write
			ack_fifo_out_csr_read                                   => mm_interconnect_0_ack_fifo_out_csr_read,                           --                                                  .read
			ack_fifo_out_csr_readdata                               => mm_interconnect_0_ack_fifo_out_csr_readdata,                       --                                                  .readdata
			ack_fifo_out_csr_writedata                              => mm_interconnect_0_ack_fifo_out_csr_writedata,                      --                                                  .writedata
			manager_debug_mem_slave_address                         => mm_interconnect_0_manager_debug_mem_slave_address,                 --                           manager_debug_mem_slave.address
			manager_debug_mem_slave_write                           => mm_interconnect_0_manager_debug_mem_slave_write,                   --                                                  .write
			manager_debug_mem_slave_read                            => mm_interconnect_0_manager_debug_mem_slave_read,                    --                                                  .read
			manager_debug_mem_slave_readdata                        => mm_interconnect_0_manager_debug_mem_slave_readdata,                --                                                  .readdata
			manager_debug_mem_slave_writedata                       => mm_interconnect_0_manager_debug_mem_slave_writedata,               --                                                  .writedata
			manager_debug_mem_slave_byteenable                      => mm_interconnect_0_manager_debug_mem_slave_byteenable,              --                                                  .byteenable
			manager_debug_mem_slave_waitrequest                     => mm_interconnect_0_manager_debug_mem_slave_waitrequest,             --                                                  .waitrequest
			manager_debug_mem_slave_debugaccess                     => mm_interconnect_0_manager_debug_mem_slave_debugaccess,             --                                                  .debugaccess
			manager_jtag_uart_avalon_jtag_slave_address             => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_address,     --               manager_jtag_uart_avalon_jtag_slave.address
			manager_jtag_uart_avalon_jtag_slave_write               => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write,       --                                                  .write
			manager_jtag_uart_avalon_jtag_slave_read                => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read,        --                                                  .read
			manager_jtag_uart_avalon_jtag_slave_readdata            => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_readdata,    --                                                  .readdata
			manager_jtag_uart_avalon_jtag_slave_writedata           => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_writedata,   --                                                  .writedata
			manager_jtag_uart_avalon_jtag_slave_waitrequest         => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_waitrequest, --                                                  .waitrequest
			manager_jtag_uart_avalon_jtag_slave_chipselect          => mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_chipselect,  --                                                  .chipselect
			mutex_s1_address                                        => mm_interconnect_0_mutex_s1_address,                                --                                          mutex_s1.address
			mutex_s1_write                                          => mm_interconnect_0_mutex_s1_write,                                  --                                                  .write
			mutex_s1_read                                           => mm_interconnect_0_mutex_s1_read,                                   --                                                  .read
			mutex_s1_readdata                                       => mm_interconnect_0_mutex_s1_readdata,                               --                                                  .readdata
			mutex_s1_writedata                                      => mm_interconnect_0_mutex_s1_writedata,                              --                                                  .writedata
			mutex_s1_chipselect                                     => mm_interconnect_0_mutex_s1_chipselect,                             --                                                  .chipselect
			pcu_control_slave_address                               => mm_interconnect_0_pcu_control_slave_address,                       --                                 pcu_control_slave.address
			pcu_control_slave_write                                 => mm_interconnect_0_pcu_control_slave_write,                         --                                                  .write
			pcu_control_slave_readdata                              => mm_interconnect_0_pcu_control_slave_readdata,                      --                                                  .readdata
			pcu_control_slave_writedata                             => mm_interconnect_0_pcu_control_slave_writedata,                     --                                                  .writedata
			pcu_control_slave_begintransfer                         => mm_interconnect_0_pcu_control_slave_begintransfer,                 --                                                  .begintransfer
			pll_0_pll_slave_address                                 => mm_interconnect_0_pll_0_pll_slave_address,                         --                                   pll_0_pll_slave.address
			pll_0_pll_slave_write                                   => mm_interconnect_0_pll_0_pll_slave_write,                           --                                                  .write
			pll_0_pll_slave_read                                    => mm_interconnect_0_pll_0_pll_slave_read,                            --                                                  .read
			pll_0_pll_slave_readdata                                => mm_interconnect_0_pll_0_pll_slave_readdata,                        --                                                  .readdata
			pll_0_pll_slave_writedata                               => mm_interconnect_0_pll_0_pll_slave_writedata,                       --                                                  .writedata
			sdram_s1_address                                        => mm_interconnect_0_sdram_s1_address,                                --                                          sdram_s1.address
			sdram_s1_write                                          => mm_interconnect_0_sdram_s1_write,                                  --                                                  .write
			sdram_s1_read                                           => mm_interconnect_0_sdram_s1_read,                                   --                                                  .read
			sdram_s1_readdata                                       => mm_interconnect_0_sdram_s1_readdata,                               --                                                  .readdata
			sdram_s1_writedata                                      => mm_interconnect_0_sdram_s1_writedata,                              --                                                  .writedata
			sdram_s1_byteenable                                     => mm_interconnect_0_sdram_s1_byteenable,                             --                                                  .byteenable
			sdram_s1_readdatavalid                                  => mm_interconnect_0_sdram_s1_readdatavalid,                          --                                                  .readdatavalid
			sdram_s1_waitrequest                                    => mm_interconnect_0_sdram_s1_waitrequest,                            --                                                  .waitrequest
			sdram_s1_chipselect                                     => mm_interconnect_0_sdram_s1_chipselect,                             --                                                  .chipselect
			shared_ocm_s1_address                                   => mm_interconnect_0_shared_ocm_s1_address,                           --                                     shared_ocm_s1.address
			shared_ocm_s1_write                                     => mm_interconnect_0_shared_ocm_s1_write,                             --                                                  .write
			shared_ocm_s1_readdata                                  => mm_interconnect_0_shared_ocm_s1_readdata,                          --                                                  .readdata
			shared_ocm_s1_writedata                                 => mm_interconnect_0_shared_ocm_s1_writedata,                         --                                                  .writedata
			shared_ocm_s1_byteenable                                => mm_interconnect_0_shared_ocm_s1_byteenable,                        --                                                  .byteenable
			shared_ocm_s1_chipselect                                => mm_interconnect_0_shared_ocm_s1_chipselect,                        --                                                  .chipselect
			shared_ocm_s1_clken                                     => mm_interconnect_0_shared_ocm_s1_clken,                             --                                                  .clken
			shared_ocm_s2_address                                   => mm_interconnect_0_shared_ocm_s2_address,                           --                                     shared_ocm_s2.address
			shared_ocm_s2_write                                     => mm_interconnect_0_shared_ocm_s2_write,                             --                                                  .write
			shared_ocm_s2_readdata                                  => mm_interconnect_0_shared_ocm_s2_readdata,                          --                                                  .readdata
			shared_ocm_s2_writedata                                 => mm_interconnect_0_shared_ocm_s2_writedata,                         --                                                  .writedata
			shared_ocm_s2_byteenable                                => mm_interconnect_0_shared_ocm_s2_byteenable,                        --                                                  .byteenable
			shared_ocm_s2_chipselect                                => mm_interconnect_0_shared_ocm_s2_chipselect,                        --                                                  .chipselect
			shared_ocm_s2_clken                                     => mm_interconnect_0_shared_ocm_s2_clken                              --                                                  .clken
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => pll_0_c0_clk,                   --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => manager_irq_irq                 --    sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => pll_0_c0_clk,                       --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of system
