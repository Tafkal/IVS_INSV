-- system_workers.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_workers is
	port (
		clk_clk            : in  std_logic                     := '0';             --   clk.clk
		reset_reset_n      : in  std_logic                     := '0';             -- reset.reset_n
		wout_waitrequest   : in  std_logic                     := '0';             --  wout.waitrequest
		wout_readdata      : in  std_logic_vector(31 downto 0) := (others => '0'); --      .readdata
		wout_readdatavalid : in  std_logic                     := '0';             --      .readdatavalid
		wout_burstcount    : out std_logic_vector(0 downto 0);                     --      .burstcount
		wout_writedata     : out std_logic_vector(31 downto 0);                    --      .writedata
		wout_address       : out std_logic_vector(27 downto 0);                    --      .address
		wout_write         : out std_logic;                                        --      .write
		wout_read          : out std_logic;                                        --      .read
		wout_byteenable    : out std_logic_vector(3 downto 0);                     --      .byteenable
		wout_debugaccess   : out std_logic                                         --      .debugaccess
	);
end entity system_workers;

architecture rtl of system_workers is
	component system_workers_cpu_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(28 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_workers_cpu_0;

	component system_workers_cpu_1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(28 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_workers_cpu_1;

	component system_workers_cpu_2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(28 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_workers_cpu_2;

	component system_workers_cpu_3 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(28 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_workers_cpu_3;

	component system_manager_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_manager_jtag_uart;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(27 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component system_workers_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			cpu_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			cpu_0_data_master_address                 : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_0_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_0_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_0_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_0_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			cpu_0_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_0_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_0_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_0_instruction_master_address          : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_0_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_0_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_0_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_address                 : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_1_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_1_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_1_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_1_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_1_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_1_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_1_instruction_master_address          : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_1_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_1_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_1_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			cpu_2_data_master_address                 : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_2_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_2_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_2_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_2_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_2_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			cpu_2_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_2_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_2_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_2_instruction_master_address          : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_2_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_2_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_2_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_2_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			cpu_3_data_master_address                 : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_3_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_3_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_3_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_3_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_3_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			cpu_3_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_3_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_3_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_3_instruction_master_address          : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			cpu_3_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_3_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_3_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_3_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			cpu_0_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_0_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_0_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_0_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_0_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_0_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_0_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_0_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			cpu_1_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_1_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_1_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_1_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_1_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_1_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_1_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_1_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			cpu_2_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_2_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_2_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_2_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_2_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_2_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_2_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_2_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			cpu_3_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_3_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_3_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_3_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_3_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_3_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_3_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_3_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			jtag_uart_0_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			jtag_uart_1_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_1_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_1_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_1_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_1_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_1_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_1_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			jtag_uart_2_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_2_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_2_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_2_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_2_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_2_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_2_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			jtag_uart_3_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_3_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_3_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_3_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_3_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_3_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_3_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			worker_out_s0_address                     : out std_logic_vector(27 downto 0);                    -- address
			worker_out_s0_write                       : out std_logic;                                        -- write
			worker_out_s0_read                        : out std_logic;                                        -- read
			worker_out_s0_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			worker_out_s0_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			worker_out_s0_burstcount                  : out std_logic_vector(0 downto 0);                     -- burstcount
			worker_out_s0_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			worker_out_s0_readdatavalid               : in  std_logic                     := 'X';             -- readdatavalid
			worker_out_s0_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			worker_out_s0_debugaccess                 : out std_logic                                         -- debugaccess
		);
	end component system_workers_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_in4      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_0_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	signal cpu_0_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	signal cpu_0_data_master_debugaccess                                   : std_logic;                     -- cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	signal cpu_0_data_master_address                                       : std_logic_vector(28 downto 0); -- cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	signal cpu_0_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	signal cpu_0_data_master_read                                          : std_logic;                     -- cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	signal cpu_0_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	signal cpu_0_data_master_write                                         : std_logic;                     -- cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	signal cpu_0_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	signal cpu_0_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	signal cpu_0_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	signal cpu_0_instruction_master_address                                : std_logic_vector(28 downto 0); -- cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	signal cpu_0_instruction_master_read                                   : std_logic;                     -- cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	signal cpu_0_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	signal cpu_3_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_3_data_master_readdata -> cpu_3:d_readdata
	signal cpu_3_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_3_data_master_waitrequest -> cpu_3:d_waitrequest
	signal cpu_3_data_master_debugaccess                                   : std_logic;                     -- cpu_3:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_3_data_master_debugaccess
	signal cpu_3_data_master_address                                       : std_logic_vector(28 downto 0); -- cpu_3:d_address -> mm_interconnect_0:cpu_3_data_master_address
	signal cpu_3_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu_3:d_byteenable -> mm_interconnect_0:cpu_3_data_master_byteenable
	signal cpu_3_data_master_read                                          : std_logic;                     -- cpu_3:d_read -> mm_interconnect_0:cpu_3_data_master_read
	signal cpu_3_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_3_data_master_readdatavalid -> cpu_3:d_readdatavalid
	signal cpu_3_data_master_write                                         : std_logic;                     -- cpu_3:d_write -> mm_interconnect_0:cpu_3_data_master_write
	signal cpu_3_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu_3:d_writedata -> mm_interconnect_0:cpu_3_data_master_writedata
	signal cpu_2_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_2_data_master_readdata -> cpu_2:d_readdata
	signal cpu_2_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_2_data_master_waitrequest -> cpu_2:d_waitrequest
	signal cpu_2_data_master_debugaccess                                   : std_logic;                     -- cpu_2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_2_data_master_debugaccess
	signal cpu_2_data_master_address                                       : std_logic_vector(28 downto 0); -- cpu_2:d_address -> mm_interconnect_0:cpu_2_data_master_address
	signal cpu_2_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu_2:d_byteenable -> mm_interconnect_0:cpu_2_data_master_byteenable
	signal cpu_2_data_master_read                                          : std_logic;                     -- cpu_2:d_read -> mm_interconnect_0:cpu_2_data_master_read
	signal cpu_2_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_2_data_master_readdatavalid -> cpu_2:d_readdatavalid
	signal cpu_2_data_master_write                                         : std_logic;                     -- cpu_2:d_write -> mm_interconnect_0:cpu_2_data_master_write
	signal cpu_2_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu_2:d_writedata -> mm_interconnect_0:cpu_2_data_master_writedata
	signal cpu_1_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	signal cpu_1_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	signal cpu_1_data_master_debugaccess                                   : std_logic;                     -- cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	signal cpu_1_data_master_address                                       : std_logic_vector(28 downto 0); -- cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	signal cpu_1_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	signal cpu_1_data_master_read                                          : std_logic;                     -- cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	signal cpu_1_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	signal cpu_1_data_master_write                                         : std_logic;                     -- cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	signal cpu_1_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	signal cpu_3_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_3_instruction_master_readdata -> cpu_3:i_readdata
	signal cpu_3_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_3_instruction_master_waitrequest -> cpu_3:i_waitrequest
	signal cpu_3_instruction_master_address                                : std_logic_vector(28 downto 0); -- cpu_3:i_address -> mm_interconnect_0:cpu_3_instruction_master_address
	signal cpu_3_instruction_master_read                                   : std_logic;                     -- cpu_3:i_read -> mm_interconnect_0:cpu_3_instruction_master_read
	signal cpu_3_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_3_instruction_master_readdatavalid -> cpu_3:i_readdatavalid
	signal cpu_2_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_2_instruction_master_readdata -> cpu_2:i_readdata
	signal cpu_2_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_2_instruction_master_waitrequest -> cpu_2:i_waitrequest
	signal cpu_2_instruction_master_address                                : std_logic_vector(28 downto 0); -- cpu_2:i_address -> mm_interconnect_0:cpu_2_instruction_master_address
	signal cpu_2_instruction_master_read                                   : std_logic;                     -- cpu_2:i_read -> mm_interconnect_0:cpu_2_instruction_master_read
	signal cpu_2_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_2_instruction_master_readdatavalid -> cpu_2:i_readdatavalid
	signal cpu_1_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	signal cpu_1_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	signal cpu_1_instruction_master_address                                : std_logic_vector(28 downto 0); -- cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	signal cpu_1_instruction_master_read                                   : std_logic;                     -- cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	signal cpu_1_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest             : std_logic;                     -- cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_0_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	signal mm_interconnect_0_cpu_0_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_0_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	signal mm_interconnect_0_cpu_0_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	signal mm_interconnect_0_worker_out_s0_readdata                        : std_logic_vector(31 downto 0); -- worker_out:s0_readdata -> mm_interconnect_0:worker_out_s0_readdata
	signal mm_interconnect_0_worker_out_s0_waitrequest                     : std_logic;                     -- worker_out:s0_waitrequest -> mm_interconnect_0:worker_out_s0_waitrequest
	signal mm_interconnect_0_worker_out_s0_debugaccess                     : std_logic;                     -- mm_interconnect_0:worker_out_s0_debugaccess -> worker_out:s0_debugaccess
	signal mm_interconnect_0_worker_out_s0_address                         : std_logic_vector(27 downto 0); -- mm_interconnect_0:worker_out_s0_address -> worker_out:s0_address
	signal mm_interconnect_0_worker_out_s0_read                            : std_logic;                     -- mm_interconnect_0:worker_out_s0_read -> worker_out:s0_read
	signal mm_interconnect_0_worker_out_s0_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:worker_out_s0_byteenable -> worker_out:s0_byteenable
	signal mm_interconnect_0_worker_out_s0_readdatavalid                   : std_logic;                     -- worker_out:s0_readdatavalid -> mm_interconnect_0:worker_out_s0_readdatavalid
	signal mm_interconnect_0_worker_out_s0_write                           : std_logic;                     -- mm_interconnect_0:worker_out_s0_write -> worker_out:s0_write
	signal mm_interconnect_0_worker_out_s0_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:worker_out_s0_writedata -> worker_out:s0_writedata
	signal mm_interconnect_0_worker_out_s0_burstcount                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:worker_out_s0_burstcount -> worker_out:s0_burstcount
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest             : std_logic;                     -- cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_1_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	signal mm_interconnect_0_cpu_1_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	signal mm_interconnect_0_cpu_1_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_1_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	signal mm_interconnect_0_cpu_1_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_chipselect -> jtag_uart_2:av_chipselect
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_2:av_readdata -> mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_2:av_waitrequest -> mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_address -> jtag_uart_2:av_address
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_writedata -> jtag_uart_2:av_writedata
	signal mm_interconnect_0_cpu_2_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu_2:debug_mem_slave_readdata -> mm_interconnect_0:cpu_2_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest             : std_logic;                     -- cpu_2:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_2_debug_mem_slave_debugaccess -> cpu_2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_2_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_2_debug_mem_slave_address -> cpu_2:debug_mem_slave_address
	signal mm_interconnect_0_cpu_2_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_2_debug_mem_slave_read -> cpu_2:debug_mem_slave_read
	signal mm_interconnect_0_cpu_2_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_2_debug_mem_slave_byteenable -> cpu_2:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_2_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_2_debug_mem_slave_write -> cpu_2:debug_mem_slave_write
	signal mm_interconnect_0_cpu_2_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_2_debug_mem_slave_writedata -> cpu_2:debug_mem_slave_writedata
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_chipselect -> jtag_uart_3:av_chipselect
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_3:av_readdata -> mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_3:av_waitrequest -> mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_address -> jtag_uart_3:av_address
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_3_avalon_jtag_slave_writedata -> jtag_uart_3:av_writedata
	signal mm_interconnect_0_cpu_3_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu_3:debug_mem_slave_readdata -> mm_interconnect_0:cpu_3_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest             : std_logic;                     -- cpu_3:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_3_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_3_debug_mem_slave_debugaccess -> cpu_3:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_3_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_3_debug_mem_slave_address -> cpu_3:debug_mem_slave_address
	signal mm_interconnect_0_cpu_3_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_3_debug_mem_slave_read -> cpu_3:debug_mem_slave_read
	signal mm_interconnect_0_cpu_3_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_3_debug_mem_slave_byteenable -> cpu_3:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_3_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_3_debug_mem_slave_write -> cpu_3:debug_mem_slave_write
	signal mm_interconnect_0_cpu_3_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_3_debug_mem_slave_writedata -> cpu_3:debug_mem_slave_writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal cpu_0_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu_0:irq
	signal irq_mapper_001_receiver0_irq                                    : std_logic;                     -- jtag_uart_1:av_irq -> irq_mapper_001:receiver0_irq
	signal cpu_1_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> cpu_1:irq
	signal irq_mapper_002_receiver0_irq                                    : std_logic;                     -- jtag_uart_2:av_irq -> irq_mapper_002:receiver0_irq
	signal cpu_2_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper_002:sender_irq -> cpu_2:irq
	signal irq_mapper_003_receiver0_irq                                    : std_logic;                     -- jtag_uart_3:av_irq -> irq_mapper_003:receiver0_irq
	signal cpu_3_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper_003:sender_irq -> cpu_3:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, worker_out:reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [cpu_0:reset_req, cpu_1:reset_req, cpu_2:reset_req, cpu_3:reset_req, rst_translator:reset_req_in]
	signal cpu_0_debug_reset_request_reset                                 : std_logic;                     -- cpu_0:debug_reset_request -> rst_controller:reset_in1
	signal cpu_1_debug_reset_request_reset                                 : std_logic;                     -- cpu_1:debug_reset_request -> rst_controller:reset_in2
	signal cpu_2_debug_reset_request_reset                                 : std_logic;                     -- cpu_2:debug_reset_request -> rst_controller:reset_in3
	signal cpu_3_debug_reset_request_reset                                 : std_logic;                     -- cpu_3:debug_reset_request -> rst_controller:reset_in4
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read:inv -> jtag_uart_1:av_read_n
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write:inv -> jtag_uart_1:av_write_n
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read:inv -> jtag_uart_2:av_read_n
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write:inv -> jtag_uart_2:av_write_n
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read:inv -> jtag_uart_3:av_read_n
	signal mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write:inv -> jtag_uart_3:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu_0:reset_n, cpu_1:reset_n, cpu_2:reset_n, cpu_3:reset_n, jtag_uart_0:rst_n, jtag_uart_1:rst_n, jtag_uart_2:rst_n, jtag_uart_3:rst_n]

begin

	cpu_0 : component system_workers_cpu_0
		port map (
			clk                                 => clk_clk,                                             --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_0_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_0_data_master_read,                              --                          .read
			d_readdata                          => cpu_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_0_data_master_write,                             --                          .write
			d_writedata                         => cpu_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_0_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_1 : component system_workers_cpu_1
		port map (
			clk                                 => clk_clk,                                             --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_1_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_1_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_1_data_master_read,                              --                          .read
			d_readdata                          => cpu_1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_1_data_master_write,                             --                          .write
			d_writedata                         => cpu_1_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_1_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_1_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_1_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_1_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_1_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_2 : component system_workers_cpu_2
		port map (
			clk                                 => clk_clk,                                             --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_2_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_2_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_2_data_master_read,                              --                          .read
			d_readdata                          => cpu_2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_2_data_master_write,                             --                          .write
			d_writedata                         => cpu_2_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_2_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_2_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_2_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_3 : component system_workers_cpu_3
		port map (
			clk                                 => clk_clk,                                             --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_3_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_3_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_3_data_master_read,                              --                          .read
			d_readdata                          => cpu_3_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_3_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_3_data_master_write,                             --                          .write
			d_writedata                         => cpu_3_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_3_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_3_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_3_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_3_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_3_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_3_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_3_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_3_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_3_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_3_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_3_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_3_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_3_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_3_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_3_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	jtag_uart_0 : component system_manager_jtag_uart
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	jtag_uart_1 : component system_manager_jtag_uart
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver0_irq                                     --               irq.irq
		);

	jtag_uart_2 : component system_manager_jtag_uart
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_002_receiver0_irq                                     --               irq.irq
		);

	jtag_uart_3 : component system_manager_jtag_uart
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_003_receiver0_irq                                     --               irq.irq
		);

	worker_out : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 28,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_clk,                                       --   clk.clk
			reset            => rst_controller_reset_out_reset,                -- reset.reset
			s0_waitrequest   => mm_interconnect_0_worker_out_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_worker_out_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_0_worker_out_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_0_worker_out_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_0_worker_out_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_0_worker_out_s0_address,       --      .address
			s0_write         => mm_interconnect_0_worker_out_s0_write,         --      .write
			s0_read          => mm_interconnect_0_worker_out_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_0_worker_out_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_0_worker_out_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => wout_waitrequest,                              --    m0.waitrequest
			m0_readdata      => wout_readdata,                                 --      .readdata
			m0_readdatavalid => wout_readdatavalid,                            --      .readdatavalid
			m0_burstcount    => wout_burstcount,                               --      .burstcount
			m0_writedata     => wout_writedata,                                --      .writedata
			m0_address       => wout_address,                                  --      .address
			m0_write         => wout_write,                                    --      .write
			m0_read          => wout_read,                                     --      .read
			m0_byteenable    => wout_byteenable,                               --      .byteenable
			m0_debugaccess   => wout_debugaccess,                              --      .debugaccess
			s0_response      => open,                                          -- (terminated)
			m0_response      => "00"                                           -- (terminated)
		);

	mm_interconnect_0 : component system_workers_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                                     --                         clk_0_clk.clk
			cpu_0_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                              -- cpu_0_reset_reset_bridge_in_reset.reset
			cpu_0_data_master_address                 => cpu_0_data_master_address,                                   --                 cpu_0_data_master.address
			cpu_0_data_master_waitrequest             => cpu_0_data_master_waitrequest,                               --                                  .waitrequest
			cpu_0_data_master_byteenable              => cpu_0_data_master_byteenable,                                --                                  .byteenable
			cpu_0_data_master_read                    => cpu_0_data_master_read,                                      --                                  .read
			cpu_0_data_master_readdata                => cpu_0_data_master_readdata,                                  --                                  .readdata
			cpu_0_data_master_readdatavalid           => cpu_0_data_master_readdatavalid,                             --                                  .readdatavalid
			cpu_0_data_master_write                   => cpu_0_data_master_write,                                     --                                  .write
			cpu_0_data_master_writedata               => cpu_0_data_master_writedata,                                 --                                  .writedata
			cpu_0_data_master_debugaccess             => cpu_0_data_master_debugaccess,                               --                                  .debugaccess
			cpu_0_instruction_master_address          => cpu_0_instruction_master_address,                            --          cpu_0_instruction_master.address
			cpu_0_instruction_master_waitrequest      => cpu_0_instruction_master_waitrequest,                        --                                  .waitrequest
			cpu_0_instruction_master_read             => cpu_0_instruction_master_read,                               --                                  .read
			cpu_0_instruction_master_readdata         => cpu_0_instruction_master_readdata,                           --                                  .readdata
			cpu_0_instruction_master_readdatavalid    => cpu_0_instruction_master_readdatavalid,                      --                                  .readdatavalid
			cpu_1_data_master_address                 => cpu_1_data_master_address,                                   --                 cpu_1_data_master.address
			cpu_1_data_master_waitrequest             => cpu_1_data_master_waitrequest,                               --                                  .waitrequest
			cpu_1_data_master_byteenable              => cpu_1_data_master_byteenable,                                --                                  .byteenable
			cpu_1_data_master_read                    => cpu_1_data_master_read,                                      --                                  .read
			cpu_1_data_master_readdata                => cpu_1_data_master_readdata,                                  --                                  .readdata
			cpu_1_data_master_readdatavalid           => cpu_1_data_master_readdatavalid,                             --                                  .readdatavalid
			cpu_1_data_master_write                   => cpu_1_data_master_write,                                     --                                  .write
			cpu_1_data_master_writedata               => cpu_1_data_master_writedata,                                 --                                  .writedata
			cpu_1_data_master_debugaccess             => cpu_1_data_master_debugaccess,                               --                                  .debugaccess
			cpu_1_instruction_master_address          => cpu_1_instruction_master_address,                            --          cpu_1_instruction_master.address
			cpu_1_instruction_master_waitrequest      => cpu_1_instruction_master_waitrequest,                        --                                  .waitrequest
			cpu_1_instruction_master_read             => cpu_1_instruction_master_read,                               --                                  .read
			cpu_1_instruction_master_readdata         => cpu_1_instruction_master_readdata,                           --                                  .readdata
			cpu_1_instruction_master_readdatavalid    => cpu_1_instruction_master_readdatavalid,                      --                                  .readdatavalid
			cpu_2_data_master_address                 => cpu_2_data_master_address,                                   --                 cpu_2_data_master.address
			cpu_2_data_master_waitrequest             => cpu_2_data_master_waitrequest,                               --                                  .waitrequest
			cpu_2_data_master_byteenable              => cpu_2_data_master_byteenable,                                --                                  .byteenable
			cpu_2_data_master_read                    => cpu_2_data_master_read,                                      --                                  .read
			cpu_2_data_master_readdata                => cpu_2_data_master_readdata,                                  --                                  .readdata
			cpu_2_data_master_readdatavalid           => cpu_2_data_master_readdatavalid,                             --                                  .readdatavalid
			cpu_2_data_master_write                   => cpu_2_data_master_write,                                     --                                  .write
			cpu_2_data_master_writedata               => cpu_2_data_master_writedata,                                 --                                  .writedata
			cpu_2_data_master_debugaccess             => cpu_2_data_master_debugaccess,                               --                                  .debugaccess
			cpu_2_instruction_master_address          => cpu_2_instruction_master_address,                            --          cpu_2_instruction_master.address
			cpu_2_instruction_master_waitrequest      => cpu_2_instruction_master_waitrequest,                        --                                  .waitrequest
			cpu_2_instruction_master_read             => cpu_2_instruction_master_read,                               --                                  .read
			cpu_2_instruction_master_readdata         => cpu_2_instruction_master_readdata,                           --                                  .readdata
			cpu_2_instruction_master_readdatavalid    => cpu_2_instruction_master_readdatavalid,                      --                                  .readdatavalid
			cpu_3_data_master_address                 => cpu_3_data_master_address,                                   --                 cpu_3_data_master.address
			cpu_3_data_master_waitrequest             => cpu_3_data_master_waitrequest,                               --                                  .waitrequest
			cpu_3_data_master_byteenable              => cpu_3_data_master_byteenable,                                --                                  .byteenable
			cpu_3_data_master_read                    => cpu_3_data_master_read,                                      --                                  .read
			cpu_3_data_master_readdata                => cpu_3_data_master_readdata,                                  --                                  .readdata
			cpu_3_data_master_readdatavalid           => cpu_3_data_master_readdatavalid,                             --                                  .readdatavalid
			cpu_3_data_master_write                   => cpu_3_data_master_write,                                     --                                  .write
			cpu_3_data_master_writedata               => cpu_3_data_master_writedata,                                 --                                  .writedata
			cpu_3_data_master_debugaccess             => cpu_3_data_master_debugaccess,                               --                                  .debugaccess
			cpu_3_instruction_master_address          => cpu_3_instruction_master_address,                            --          cpu_3_instruction_master.address
			cpu_3_instruction_master_waitrequest      => cpu_3_instruction_master_waitrequest,                        --                                  .waitrequest
			cpu_3_instruction_master_read             => cpu_3_instruction_master_read,                               --                                  .read
			cpu_3_instruction_master_readdata         => cpu_3_instruction_master_readdata,                           --                                  .readdata
			cpu_3_instruction_master_readdatavalid    => cpu_3_instruction_master_readdatavalid,                      --                                  .readdatavalid
			cpu_0_debug_mem_slave_address             => mm_interconnect_0_cpu_0_debug_mem_slave_address,             --             cpu_0_debug_mem_slave.address
			cpu_0_debug_mem_slave_write               => mm_interconnect_0_cpu_0_debug_mem_slave_write,               --                                  .write
			cpu_0_debug_mem_slave_read                => mm_interconnect_0_cpu_0_debug_mem_slave_read,                --                                  .read
			cpu_0_debug_mem_slave_readdata            => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,            --                                  .readdata
			cpu_0_debug_mem_slave_writedata           => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,           --                                  .writedata
			cpu_0_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,          --                                  .byteenable
			cpu_0_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest,         --                                  .waitrequest
			cpu_0_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess,         --                                  .debugaccess
			cpu_1_debug_mem_slave_address             => mm_interconnect_0_cpu_1_debug_mem_slave_address,             --             cpu_1_debug_mem_slave.address
			cpu_1_debug_mem_slave_write               => mm_interconnect_0_cpu_1_debug_mem_slave_write,               --                                  .write
			cpu_1_debug_mem_slave_read                => mm_interconnect_0_cpu_1_debug_mem_slave_read,                --                                  .read
			cpu_1_debug_mem_slave_readdata            => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,            --                                  .readdata
			cpu_1_debug_mem_slave_writedata           => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,           --                                  .writedata
			cpu_1_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,          --                                  .byteenable
			cpu_1_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest,         --                                  .waitrequest
			cpu_1_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess,         --                                  .debugaccess
			cpu_2_debug_mem_slave_address             => mm_interconnect_0_cpu_2_debug_mem_slave_address,             --             cpu_2_debug_mem_slave.address
			cpu_2_debug_mem_slave_write               => mm_interconnect_0_cpu_2_debug_mem_slave_write,               --                                  .write
			cpu_2_debug_mem_slave_read                => mm_interconnect_0_cpu_2_debug_mem_slave_read,                --                                  .read
			cpu_2_debug_mem_slave_readdata            => mm_interconnect_0_cpu_2_debug_mem_slave_readdata,            --                                  .readdata
			cpu_2_debug_mem_slave_writedata           => mm_interconnect_0_cpu_2_debug_mem_slave_writedata,           --                                  .writedata
			cpu_2_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_2_debug_mem_slave_byteenable,          --                                  .byteenable
			cpu_2_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest,         --                                  .waitrequest
			cpu_2_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess,         --                                  .debugaccess
			cpu_3_debug_mem_slave_address             => mm_interconnect_0_cpu_3_debug_mem_slave_address,             --             cpu_3_debug_mem_slave.address
			cpu_3_debug_mem_slave_write               => mm_interconnect_0_cpu_3_debug_mem_slave_write,               --                                  .write
			cpu_3_debug_mem_slave_read                => mm_interconnect_0_cpu_3_debug_mem_slave_read,                --                                  .read
			cpu_3_debug_mem_slave_readdata            => mm_interconnect_0_cpu_3_debug_mem_slave_readdata,            --                                  .readdata
			cpu_3_debug_mem_slave_writedata           => mm_interconnect_0_cpu_3_debug_mem_slave_writedata,           --                                  .writedata
			cpu_3_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_3_debug_mem_slave_byteenable,          --                                  .byteenable
			cpu_3_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest,         --                                  .waitrequest
			cpu_3_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess,         --                                  .debugaccess
			jtag_uart_0_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --     jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_0_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_0_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_0_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                  .chipselect
			jtag_uart_1_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address,     --     jtag_uart_1_avalon_jtag_slave.address
			jtag_uart_1_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_1_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_1_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_1_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_1_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_1_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect,  --                                  .chipselect
			jtag_uart_2_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_address,     --     jtag_uart_2_avalon_jtag_slave.address
			jtag_uart_2_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_2_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_2_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_2_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_2_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_2_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_chipselect,  --                                  .chipselect
			jtag_uart_3_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_address,     --     jtag_uart_3_avalon_jtag_slave.address
			jtag_uart_3_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_3_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_3_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_3_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_3_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_3_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_chipselect,  --                                  .chipselect
			worker_out_s0_address                     => mm_interconnect_0_worker_out_s0_address,                     --                     worker_out_s0.address
			worker_out_s0_write                       => mm_interconnect_0_worker_out_s0_write,                       --                                  .write
			worker_out_s0_read                        => mm_interconnect_0_worker_out_s0_read,                        --                                  .read
			worker_out_s0_readdata                    => mm_interconnect_0_worker_out_s0_readdata,                    --                                  .readdata
			worker_out_s0_writedata                   => mm_interconnect_0_worker_out_s0_writedata,                   --                                  .writedata
			worker_out_s0_burstcount                  => mm_interconnect_0_worker_out_s0_burstcount,                  --                                  .burstcount
			worker_out_s0_byteenable                  => mm_interconnect_0_worker_out_s0_byteenable,                  --                                  .byteenable
			worker_out_s0_readdatavalid               => mm_interconnect_0_worker_out_s0_readdatavalid,               --                                  .readdatavalid
			worker_out_s0_waitrequest                 => mm_interconnect_0_worker_out_s0_waitrequest,                 --                                  .waitrequest
			worker_out_s0_debugaccess                 => mm_interconnect_0_worker_out_s0_debugaccess                  --                                  .debugaccess
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => cpu_0_irq_irq                   --    sender.irq
		);

	irq_mapper_001 : component system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,   -- receiver0.irq
			sender_irq    => cpu_1_irq_irq                   --    sender.irq
		);

	irq_mapper_002 : component system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_002_receiver0_irq,   -- receiver0.irq
			sender_irq    => cpu_2_irq_irq                   --    sender.irq
		);

	irq_mapper_003 : component system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_003_receiver0_irq,   -- receiver0.irq
			sender_irq    => cpu_3_irq_irq                   --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 5,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_0_debug_reset_request_reset,    -- reset_in1.reset
			reset_in2      => cpu_1_debug_reset_request_reset,    -- reset_in2.reset
			reset_in3      => cpu_2_debug_reset_request_reset,    -- reset_in3.reset
			reset_in4      => cpu_3_debug_reset_request_reset,    -- reset_in4.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_3_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of system_workers
